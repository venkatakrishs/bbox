/****** Imports *******/
import bbox_types :: *;

/*********************/


function BBoxOutput fn_compute(BBoxInput inp);
  BBoxOutput result = unpack(0);
  return result;
endfunction
